//-----------------------------------------------------------------------------
//
// Title       : IULogical
// Design      : SPARC
// Author      : Dina
// Company     : Dina
//
//-----------------------------------------------------------------------------
//
// File        : IULogical.v
// Generated   : Thu Jun 13 02:59:02 2013
// From        : interface description file
// By          : Itf2Vhdl ver. 1.22
//
//-----------------------------------------------------------------------------
//
// Description : 
//
//-----------------------------------------------------------------------------
`timescale 1 ns / 1 ps

//{{ Section below this comment is automatically maintained
//   and may be overwritten
//{module {IULogical}}
module IULogical ();
//}} End of automatically maintained section

// -- Enter your statements here -- //

endmodule
